$date
	Fri Jul 31 20:20:15 2020
$end
$version
	Icarus Verilog
$end
$timescale
	1ps
$end
$scope module Tabla1POS $end
$var wire 1 ! NA $end
$var wire 1 " NB $end
$var wire 1 # NC $end
$var wire 1 $ P1 $end
$var wire 1 % S1 $end
$var wire 1 & S2 $end
$var wire 1 ' S3 $end
$var reg 1 ( A $end
$var reg 1 ) B $end
$var reg 1 * C $end
$upscope $end
$enddefinitions $end
#0
$dumpvars
0*
0)
0(
1'
1&
1%
1$
1#
1"
1!
$end
#1
0$
0%
0#
1*
#2
1$
1#
1%
0"
0*
1)
#3
0$
0&
0#
1*
#4
1$
1#
1"
1&
0!
0*
0)
1(
#5
0#
1*
#6
0$
0'
1#
0"
0*
1)
#7
1$
1'
0#
1*
#8
